-- Copyright (C) 1991-2010 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 9.1 Build 304 01/25/2010 Service Pack 1 SJ Web Edition
-- Created on Fri Aug 13 13:08:55 2021

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY collis IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        w : IN STD_LOGIC := '0';
        z : OUT STD_LOGIC
    );
END collis;

ARCHITECTURE BEHAVIOR OF collis IS
    TYPE type_fstate IS (s0,s1,s2,s3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,w)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= s0;
            z <= '0';
        ELSE
            z <= '0';
            CASE fstate IS
                WHEN s0 =>
                    IF (NOT((w = '1'))) THEN
                        reg_fstate <= s0;
                    ELSIF ((w = '1')) THEN
                        reg_fstate <= s1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= s0;
                    END IF;

                    IF (NOT((w = '1'))) THEN
                        z <= '0';
                    ELSIF ((w = '1')) THEN
                        z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z <= '0';
                    END IF;
                WHEN s1 =>
                    IF ((w = '1')) THEN
                        reg_fstate <= s2;
                    ELSIF (NOT((w = '1'))) THEN
                        reg_fstate <= s3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= s1;
                    END IF;

                    IF (NOT((w = '1'))) THEN
                        z <= '0';
                    ELSIF ((w = '1')) THEN
                        z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z <= '0';
                    END IF;
                WHEN s2 =>
                    IF ((w = '1')) THEN
                        reg_fstate <= s1;
                    ELSIF (NOT((w = '1'))) THEN
                        reg_fstate <= s3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= s2;
                    END IF;

                    IF (NOT((w = '1'))) THEN
                        z <= '0';
                    ELSIF ((w = '1')) THEN
                        z <= '0';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z <= '0';
                    END IF;
                WHEN s3 =>
                    IF ((w = '1')) THEN
                        reg_fstate <= s2;
                    ELSIF (NOT((w = '1'))) THEN
                        reg_fstate <= s0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= s3;
                    END IF;

                    IF (NOT((w = '1'))) THEN
                        z <= '0';
                    ELSIF ((w = '1')) THEN
                        z <= '1';
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        z <= '0';
                    END IF;
                WHEN OTHERS => 
                    z <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
